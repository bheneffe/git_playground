UART baud_rate = 115200;
