module uart (
    input logic clk,
    input logic rst_n,
    input logic rx,
    output logic tx
);
    // UART implementation here
endmodule
