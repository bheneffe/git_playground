UART baud_rate = 9600;
